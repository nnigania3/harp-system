// Copyright (C) 1991-2012 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 12.1 Build 177 11/07/2012 SJ Web Edition
// Created on Thu Mar 14 15:27:03 2013

// synthesis message_off 10175

`timescale 1ns/1ns

module blocking (
    reset,clock,dirty,rw_prev,stall_l2,done_l2,miss,
    rw_l2,valid_l2,we_b,rd_valid_b,l2_addr_en,stall_proc);

    input reset;
    input clock;
    input dirty;
    input rw_prev;
    input stall_l2;
    input done_l2;
    input miss;
    tri0 reset;
    tri0 dirty;
    tri0 rw_prev;
    tri0 stall_l2;
    tri0 done_l2;
    tri0 miss;
    output rw_l2;
    output valid_l2;
    output we_b;
    output rd_valid_b;
    output l2_addr_en;
    output stall_proc;
    reg rw_l2;
    reg reg_rw_l2;
    reg valid_l2;
    reg reg_valid_l2;
    reg we_b;
    reg reg_we_b;
    reg rd_valid_b;
    reg reg_rd_valid_b;
    reg l2_addr_en;
    reg reg_l2_addr_en;
    reg stall_proc;
    reg reg_stall_proc;
    reg [5:0] fstate;
    reg [5:0] reg_fstate;
    parameter Idle=0,Read_l2=1,WB_L2=2,Read_L1=3,Write_L1=4,Read_Wait=5;

    initial
    begin
        reg_rw_l2 <= 1'b0;
        reg_valid_l2 <= 1'b0;
        reg_we_b <= 1'b0;
        reg_rd_valid_b <= 1'b0;
        reg_l2_addr_en <= 1'b0;
        reg_stall_proc <= 1'b0;
    end

    always @(posedge clock or negedge reset)
    begin
        if (~reset) begin
            fstate <= Idle;
            rw_l2 <= 1'b0;
            valid_l2 <= 1'b0;
            we_b <= 1'b0;
            rd_valid_b <= 1'b0;
            l2_addr_en <= 1'b0;
            stall_proc <= 1'b0;
        end
        else begin
            fstate <= reg_fstate;
            rw_l2 <= reg_rw_l2;
            valid_l2 <= reg_valid_l2;
            we_b <= reg_we_b;
            rd_valid_b <= reg_rd_valid_b;
            l2_addr_en <= reg_l2_addr_en;
            stall_proc <= reg_stall_proc;
        end
    end

    always @(fstate or dirty or rw_prev or stall_l2 or done_l2 or miss)
    begin
        reg_rw_l2 <= 1'b0;
        reg_valid_l2 <= 1'b0;
        reg_we_b <= 1'b0;
        reg_rd_valid_b <= 1'b0;
        reg_l2_addr_en <= 1'b0;
        reg_stall_proc <= 1'b0;
        case (fstate)
            Idle: begin
                if (((miss & dirty) & ~(stall_l2)))
                    reg_fstate <= WB_L2;
                else if (((miss & ~(dirty)) & ~(stall_l2)))
                    reg_fstate <= Read_l2;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= Idle;

                reg_rd_valid_b <= 1'b0;

                reg_stall_proc <= 1'b0;

                reg_we_b <= 1'b0;

                reg_valid_l2 <= 1'b0;

                reg_l2_addr_en <= 1'b0;

                reg_rw_l2 <= 1'b0;
            end
            Read_l2: begin
                reg_fstate <= Read_Wait;

                reg_stall_proc <= 1'b0;

                reg_we_b <= 1'b0;

                reg_valid_l2 <= 1'b1;

                reg_l2_addr_en <= 1'b0;

                reg_rw_l2 <= 1'b0;
            end
            WB_L2: begin
                reg_fstate <= Read_l2;

                reg_rd_valid_b <= 1'b1;

                reg_stall_proc <= 1'b0;

                reg_we_b <= 1'b0;

                reg_valid_l2 <= 1'b1;

                reg_l2_addr_en <= 1'b1;

                reg_rw_l2 <= 1'b1;
            end
            Read_L1: begin
                reg_fstate <= Idle;

                reg_stall_proc <= 1'b1;

                reg_we_b <= 1'b0;

                reg_valid_l2 <= 1'b0;
            end
            Write_L1: begin
                reg_fstate <= Idle;

                reg_stall_proc <= 1'b1;

                reg_we_b <= 1'b1;

                reg_valid_l2 <= 1'b0;
            end
            Read_Wait: begin
                if ((done_l2 & ~(rw_prev)))
                    reg_fstate <= Read_L1;
                else if ((done_l2 & rw_prev))
                    reg_fstate <= Write_L1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= Read_Wait;

                reg_stall_proc <= 1'b0;

                reg_we_b <= 1'b0;

                reg_valid_l2 <= 1'b0;
            end
            default: begin
                reg_rw_l2 <= 1'bx;
                reg_valid_l2 <= 1'bx;
                reg_we_b <= 1'bx;
                reg_rd_valid_b <= 1'bx;
                reg_l2_addr_en <= 1'bx;
                reg_stall_proc <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // blocking
